CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 120 30 200 10
1200 75 2302 1003
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 1
21 1Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1368 171 1481 268
77070354 0
0
2 

2 

0
0
0
60
13 OV7660FSL CON
94 1033 368 0 24 49
0 29 28 27 26 25 24 23 22 21
20 19 18 17 16 15 14 13 12 11
10 9 8 7 6
13 OV7660FSL CON
1 0 4992 512
12 54550-2494-C
-35 130 49 138
4 CON5
-10 -127 18 -119
33 Molex ZIF Connector for OV7660FSL
-108 -147 123 -139
0
0
0
0
13 MOLEX05FPC-24
49

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 0
0 0 0 0 1 0 0 0
3 CON
5130 0 0
2
5.89415e-315 0
0
13 OV7660FSL CON
94 1147 368 0 24 49
0 29 28 27 26 25 24 23 22 21
20 19 18 17 16 15 14 13 12 11
10 9 8 7 6
13 OV7660FSL CON
2 0 4992 0
12 54550-2494-C
-32 129 52 137
4 CON6
-4 -127 24 -119
33 Molex ZIF Connector for OV7660FSL
-108 -147 123 -139
0
0
0
0
13 MOLEX05FPC-24
49

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 0
0 0 0 0 1 0 0 0
3 CON
391 0 0
2
5.89415e-315 5.26354e-315
0
9 Terminal~
194 878 343 0 1 3
0 2
0
0 0 49504 90
4 DVdd
-32 -6 -4 2
3 T12
-11 -32 10 -24
0
5 DVdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3124 0 0
2
40299 0
0
9 Terminal~
194 702 49 0 1 3
0 2
0
0 0 49504 270
4 DVdd
-14 -15 14 -7
3 T11
-11 -32 10 -24
0
5 DVdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3421 0 0
2
40299 1
0
9 Terminal~
194 838 203 0 1 3
0 3
0
0 0 49504 0
4 AVdd
-14 -13 14 -5
3 T10
-11 -32 10 -24
0
5 AVdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8157 0 0
2
40299 2
0
9 Terminal~
194 645 40 0 1 3
0 3
0
0 0 49504 270
4 AVdd
-14 -15 14 -7
2 T9
-7 -32 7 -24
0
5 AVdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5572 0 0
2
40299 3
0
9 Terminal~
194 782 204 0 1 3
0 4
0
0 0 49504 0
3 Vdd
-11 -14 10 -6
2 T8
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8901 0 0
2
40299 4
0
9 Terminal~
194 664 516 0 1 3
0 4
0
0 0 49504 0
3 Vdd
-11 -15 10 -7
2 T7
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7361 0 0
2
40299 5
0
9 Terminal~
194 558 514 0 1 3
0 4
0
0 0 49504 90
3 Vdd
-9 -15 12 -7
2 T6
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4747 0 0
2
40299 6
0
9 Terminal~
194 191 281 0 1 3
0 4
0
0 0 49504 0
3 Vdd
-10 -15 11 -7
2 T5
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
972 0 0
2
40299 7
0
9 Terminal~
194 421 482 0 1 3
0 4
0
0 0 49504 270
3 Vdd
-19 -13 2 -5
2 T4
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3472 0 0
2
40299 8
0
9 Terminal~
194 518 369 0 1 3
0 4
0
0 0 49504 270
3 Vdd
2 -5 23 3
2 T3
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9998 0 0
2
40299 9
0
9 Terminal~
194 382 139 0 1 3
0 4
0
0 0 49504 0
3 Vdd
-10 -15 11 -7
2 T2
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3536 0 0
2
40299 10
0
9 Terminal~
194 385 52 0 1 3
0 4
0
0 0 49504 270
3 Vdd
-11 -15 10 -7
2 T1
-8 -32 6 -24
0
4 Vdd;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4597 0 0
2
40299 11
0
10 Capacitor~
219 436 143 0 2 5
0 5 64
0
0 0 832 180
5 2.2uF
-18 -18 17 -10
2 C8
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3835 0 0
2
5.89415e-315 5.30499e-315
0
7 Ground~
168 465 150 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
5.89415e-315 5.32571e-315
0
7 Ground~
168 611 89 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
40299 12
0
10 Capacitor~
219 611 66 0 2 5
0 5 3
0
0 0 832 90
3 1uF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9323 0 0
2
40299 13
0
10 Capacitor~
219 448 59 0 2 5
0 5 34
0
0 0 832 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
317 0 0
2
40299 14
0
7 Ground~
168 448 92 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
40299 15
0
10 Capacitor~
219 659 66 0 2 5
0 5 2
0
0 0 832 90
3 1uF
11 0 32 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4299 0 0
2
40299 16
0
6 SIP10~
219 153 525 0 10 21
0 5 34 47 41 40 39 38 30 37
36
0
0 0 864 782
5 Extra
-16 12 19 20
4 CON4
44 0 72 8
0
0
0
0
0
11 SIP10/SM575
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
0 0 0 0 1 0 0 0
3 CON
9672 0 0
2
5.89415e-315 5.34643e-315
0
7 Ground~
168 641 520 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
40299 17
0
5 SIP3~
219 597 451 0 3 7
0 44 45 31
0
0 0 992 0
10 OSC Source
12 -4 82 4
2 J1
-4 -25 10 -17
0
0
0
0
0
12 SM/JP/0402-3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
6369 0 0
2
40299 18
0
7 Ground~
168 816 467 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
40299 19
0
7 Ground~
168 240 424 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7100 0 0
2
40299 20
0
7 Ground~
168 369 513 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
40299 21
0
7 Ground~
168 585 349 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
40299 22
0
5 SIP5~
219 436 510 0 5 11
0 63 62 61 60 5
0
0 0 864 270
4 UART
-13 12 15 20
4 CON2
24 0 52 8
0
0
0
0
0
4 pad5
11

0 1 2 3 4 5 1 2 3 4
5 0
0 0 0 0 1 0 0 0
1 J
961 0 0
2
40299 23
0
10 Capacitor~
219 884 249 0 2 5
0 5 3
0
0 0 832 90
5 0.1uF
-42 1 -7 9
2 C6
-32 -9 -18 -1
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3178 0 0
2
40299 24
0
5 SIP5~
219 337 587 0 5 11
0 33 4 5 58 59
0
0 0 864 270
4 ICD2
-15 12 13 20
4 CON3
-53 0 -25 8
0
0
0
0
0
4 pad5
11

0 1 2 3 4 5 1 2 3 4
5 0
0 0 0 0 1 0 0 0
1 J
3409 0 0
2
40299 25
0
7 Ground~
168 95 544 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3951 0 0
2
40299 26
0
4 LED~
171 333 177 0 2 2
12 53 55
0
0 0 736 270
4 LED1
26 -14 54 -6
2 D1
9 -14 23 -6
0
0
11 %D %1 %2 %M
0
0
12 SM/D/0402/12
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8885 0 0
2
40299 27
0
4 LED~
171 334 207 0 2 2
10 52 54
0
0 0 608 270
4 LED1
-12 -20 16 -12
2 D2
10 -13 24 -5
0
0
11 %D %1 %2 %M
0
0
12 SM/D/0402/12
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3780 0 0
2
40299 28
0
7 Ground~
168 281 213 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
40299 29
0
14 NO PushButton~
191 709 606 0 2 5
0 51 5
0
0 0 4704 512
9 B3U-3100P
-31 -20 32 -12
2 S1
7 -13 21 -5
28 Side-actuated Tactile Switch
-98 -40 98 -32
0
0
0
0
9 B3U-3100P
5

0 1 2 1 2 0
0 0 0 0 1 0 -1 0
1 S
9442 0 0
2
40299 30
0
7 Ground~
168 735 632 0 1 3
0 5
0
0 0 53344 512
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9424 0 0
2
40299 31
0
14 NO PushButton~
191 709 578 0 2 5
0 50 5
0
0 0 4704 512
9 B3U-3100P
-31 -20 32 -12
2 S2
6 -15 20 -7
28 Side-actuated Tactile Switch
-98 -40 98 -32
0
0
0
0
9 B3U-3100P
5

0 1 2 1 2 0
0 0 0 0 1 0 -1 0
1 S
9968 0 0
2
40299 32
0
10 Capacitor~
219 219 390 0 2 5
0 5 4
0
0 0 832 180
5 0.1uF
-17 14 18 22
2 C7
-6 25 8 33
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9281 0 0
2
40299 33
0
10 Capacitor~
219 357 74 0 2 5
0 5 4
0
0 0 832 90
5 2.2uF
10 1 45 9
2 C5
19 -11 33 -3
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8464 0 0
2
5.89415e-315 5.3568e-315
0
7 Ground~
168 357 94 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
5.89415e-315 5.36716e-315
0
7 Ground~
168 221 96 0 1 3
0 5
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.89415e-315 5.37752e-315
0
5 SIP2~
219 37 55 0 2 5
0 5 34
0
0 0 864 180
5 ~3.7V
-26 -20 9 -12
7 BATTERY
-31 -32 18 -24
0
0
0
0
0
4 pad2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
4139 0 0
2
5.89415e-315 5.38788e-315
0
10 Capacitor~
219 221 68 0 2 5
0 5 34
0
0 0 832 90
3 1uF
11 0 32 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6435 0 0
2
5.89415e-315 5.39306e-315
0
12 ZXCL Series~
94 301 63 0 5 11
0 34 5 34 77 4
12 ZXCL Series~
3 0 4864 0
11 ZXCL330H5TA
-31 33 46 41
4 REG1
-7 -34 21 -26
38 Micropower 150mA Low-Dropout Regulator
-125 -64 141 -56
0
0
0
0
6 SC70-5
11

0 1 2 3 4 5 1 2 3 4
5 0
0 0 0 512 1 0 0 0
3 REG
5283 0 0
2
5.89415e-315 5.39824e-315
0
14 MN1380 Series~
94 150 96 0 3 7
0 35 5 34
14 MN1380 Series~
4 0 4864 180
9 MN13822-L
-43 28 20 36
4 SUP1
-27 -28 1 -20
27 Voltage Detector/Supervisor
-109 -48 80 -40
0
0
0
0
8 SC59/132
7

0 1 3 2 1 3 2 0
0 0 0 0 1 1 0 0
3 SUP
6874 0 0
2
5.89415e-315 5.40342e-315
0
13 dsPIC33FJ...~
94 390 341 0 64 129
0 78 79 80 68 65 66 33 67 5
4 81 82 41 40 39 38 59 58 4
5 60 83 84 85 5 4 86 87 61
88 62 63 48 49 35 30 37 4 31
44 5 57 56 46 36 76 42 32 75
74 73 72 71 70 69 64 53 52 89
90 47 91 92 4
13 dsPIC33FJ...~
5 0 4864 0
15 dsPIC33FJ128...
-59 -2 46 6
5 PROC1
68 -109 103 -101
17 dsPIC33FJ128MC706
-64 -132 55 -124
0
0
0
0
9 Q.50M_64A
129

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 58 59 60
61 62 63 64 57 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 58 59 60 61 62 63 64 57 0
0 0 0 512 1 0 0 0
4 PROC
5305 0 0
2
40299 34
0
11 AT45DB161D~
94 142 377 0 8 17
0 66 68 4 67 4 4 5 65
11 AT45DB161D~
6 0 4864 0
13 AT45DB161D-MU
-42 30 49 38
4 MEM1
-14 -28 14 -20
23 16Mbit DataFlash Memory
-80 -57 81 -49
0
0
0
0
5 MLF-8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
3 MEM
34 0 0
2
5.89415e-315 5.4086e-315
0
14 MIC5320 Serie~
94 540 48 0 6 13
0 34 5 32 32 2 3
13 MIC5320 Serie
7 0 4864 0
13 MIC5320-JGYML
-39 20 52 28
4 REG2
-13 -28 15 -20
37 High Performance Dual 150mA uCap ULDO
-129 -48 130 -40
0
0
0
0
5 MLF-6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 0 1 0 0 0
3 REG
969 0 0
2
5.89415e-315 5.41378e-315
0
13 OV7660FSL CON
94 910 368 0 24 49
0 93 5 30 3 37 5 57 42 56
2 3 69 45 70 5 71 46 72 76
73 75 74 94 95
13 OV7660FSL CON
8 0 4992 0
12 54550-2494-C
-25 128 59 136
4 CON1
-4 -127 24 -119
33 Molex ZIF Connector for OV7660FSL
-108 -147 123 -139
0
0
0
0
13 MOLEX05FPC-24
49

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 0
0 0 0 512 1 0 0 0
3 CON
8402 0 0
2
5.89415e-315 5.41896e-315
0
14 ECS3963 Serie~
94 611 502 0 4 9
0 96 5 31 4
14 ECS3963 Serie~
9 0 4608 180
15 ECS-3963-400-BN
-59 -19 46 -11
4 OSC1
-21 -19 7 -11
24 ECS SMD Clock Oscillator
-84 -48 84 -40
0
0
0
0
11 ECS3963_SMD
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 OSC
3751 0 0
2
5.89415e-315 5.42414e-315
0
9 Resistor~
219 764 244 0 2 5
0 30 4
0
0 0 864 90
4 4.7k
2 0 30 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4292 0 0
2
40299 35
0
9 Resistor~
219 801 243 0 2 5
0 37 4
0
0 0 864 90
4 4.7k
2 0 30 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6118 0 0
2
40299 36
0
9 Resistor~
219 385 553 0 2 5
0 33 4
0
0 0 864 90
3 10k
7 0 28 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
40299 37
0
9 Resistor~
219 308 175 0 3 5
0 5 55 -1
0
0 0 864 0
3 470
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6357 0 0
2
40299 38
0
9 Resistor~
219 308 205 0 3 5
0 5 54 -1
0
0 0 864 0
3 470
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
319 0 0
2
40299 39
0
9 Resistor~
219 616 586 0 2 5
0 49 50
0
0 0 864 0
3 470
-11 -14 10 -6
2 R7
-25 -20 -11 -12
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3976 0 0
2
40299 40
0
9 Resistor~
219 618 614 0 2 5
0 48 51
0
0 0 864 0
3 470
-11 -14 10 -6
2 R9
-28 -19 -14 -11
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7634 0 0
2
40299 41
0
9 Resistor~
219 672 559 0 2 5
0 51 4
0
0 0 864 90
3 10k
5 1 26 9
3 R10
5 -9 26 -1
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
523 0 0
2
40299 42
0
9 Resistor~
219 656 558 0 2 5
0 50 4
0
0 0 864 90
3 10k
-24 2 -3 10
2 R8
-20 -8 -6 0
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6748 0 0
2
40299 43
0
140
4 1 4 0 0 4096 0 51 9 0 0 2
574 512
569 512
24 24 6 0 0 4224 0 2 1 0 0 2
1132 467
1062 467
23 23 7 0 0 4224 0 2 1 0 0 2
1132 458
1062 458
22 22 8 0 0 4224 0 2 1 0 0 2
1132 449
1062 449
21 21 9 0 0 4224 0 2 1 0 0 2
1132 440
1062 440
20 20 10 0 0 4224 0 2 1 0 0 2
1132 431
1062 431
19 19 11 0 0 4224 0 2 1 0 0 2
1132 422
1062 422
18 18 12 0 0 4224 0 2 1 0 0 2
1132 413
1062 413
17 17 13 0 0 4224 0 2 1 0 0 2
1132 404
1062 404
16 16 14 0 0 4224 0 2 1 0 0 2
1132 395
1062 395
15 15 15 0 0 4224 0 2 1 0 0 2
1132 386
1062 386
14 14 16 0 0 4224 0 2 1 0 0 2
1132 377
1062 377
13 13 17 0 0 4224 0 2 1 0 0 2
1132 368
1062 368
12 12 18 0 0 4224 0 2 1 0 0 2
1132 359
1062 359
11 11 19 0 0 4224 0 2 1 0 0 2
1132 350
1062 350
10 10 20 0 0 4224 0 2 1 0 0 2
1132 341
1062 341
9 9 21 0 0 4224 0 2 1 0 0 2
1132 332
1062 332
8 8 22 0 0 4224 0 2 1 0 0 2
1132 323
1062 323
7 7 23 0 0 4224 0 2 1 0 0 2
1132 314
1062 314
6 6 24 0 0 4224 0 2 1 0 0 2
1132 305
1062 305
5 5 25 0 0 4224 0 2 1 0 0 2
1132 296
1062 296
4 4 26 0 0 4224 0 2 1 0 0 2
1132 287
1062 287
3 3 27 0 0 4224 0 2 1 0 0 2
1132 278
1062 278
2 2 28 0 0 4224 0 2 1 0 0 2
1132 269
1062 269
1 1 29 0 0 4224 0 2 1 0 0 2
1132 260
1062 260
1 38 4 0 0 4096 0 12 47 0 0 2
506 368
492 368
0 36 30 0 0 4096 0 0 47 122 0 2
505 386
492 386
1 0 4 0 0 0 0 7 0 0 119 2
782 213
782 216
1 2 5 0 0 4096 0 23 51 0 0 3
641 514
641 503
631 503
3 0 31 0 0 4096 0 51 0 0 68 2
574 503
574 460
6 0 5 0 0 4096 0 50 0 0 112 2
895 305
816 305
48 0 32 0 0 8320 0 47 0 0 34 3
492 278
544 278
544 84
1 1 5 0 0 0 0 16 15 0 0 3
465 144
465 143
445 143
3 4 32 0 0 0 0 49 49 0 0 6
507 57
492 57
492 84
592 84
592 57
579 57
2 0 5 0 0 0 0 49 0 0 52 4
507 48
484 48
484 78
448 78
3 0 4 0 0 12416 0 48 0 0 38 4
100 386
83 386
83 297
191 297
10 0 4 0 0 0 0 47 0 0 38 2
280 359
191 359
0 1 4 0 0 0 0 0 10 39 0 2
191 390
191 290
2 0 4 0 0 0 0 39 0 0 111 2
210 390
191 390
7 1 33 0 0 8320 0 47 31 0 0 7
280 332
278 332
278 614
385 614
385 578
354 578
354 579
1 0 5 0 0 0 0 39 0 0 42 2
228 390
240 390
9 1 5 0 0 0 0 47 26 0 0 3
280 350
240 350
240 418
0 0 34 0 0 8192 0 0 0 44 49 4
91 52
91 15
448 15
448 39
3 0 34 0 0 0 0 46 0 0 138 3
117 99
91 99
91 52
2 0 2 0 0 4096 0 21 0 0 47 2
659 57
659 48
2 0 3 0 0 4096 0 18 0 0 48 2
611 57
611 39
5 1 2 0 0 4224 0 49 4 0 0 2
579 48
690 48
6 1 3 0 0 4096 0 49 6 0 0 2
579 39
633 39
2 1 34 0 0 0 0 19 49 0 0 3
448 50
448 39
507 39
1 1 5 0 0 0 0 21 17 0 0 4
659 75
659 82
611 82
611 83
1 1 5 0 0 0 0 18 17 0 0 4
611 75
611 85
611 85
611 83
1 1 5 0 0 0 0 20 19 0 0 2
448 86
448 68
0 2 5 0 0 0 0 0 46 55 0 2
196 87
155 87
1 35 35 0 0 4224 0 46 47 0 0 4
155 111
501 111
501 395
492 395
1 0 5 0 0 4224 0 43 0 0 139 4
41 61
196 61
196 87
222 87
10 45 36 0 0 20608 0 22 47 0 0 7
190 517
190 510
237 510
237 637
542 637
542 305
492 305
9 0 37 0 0 16384 0 22 0 0 123 6
181 517
181 504
243 504
243 629
514 629
514 377
16 7 38 0 0 12416 0 47 22 0 0 5
280 413
272 413
272 490
163 490
163 517
15 6 39 0 0 12416 0 47 22 0 0 5
280 404
267 404
267 483
154 483
154 517
14 5 40 0 0 12416 0 47 22 0 0 5
280 395
261 395
261 474
145 474
145 517
13 4 41 0 0 12416 0 47 22 0 0 5
280 386
255 386
255 465
136 465
136 517
1 1 5 0 0 0 0 22 32 0 0 4
109 517
109 515
95 515
95 538
8 47 42 0 0 4224 0 50 47 0 0 4
895 323
637 323
637 287
492 287
0 2 34 0 0 4224 0 0 22 138 0 4
51 52
51 506
118 506
118 517
0 0 43 0 0 0 0 0 0 0 0 2
630 456
630 456
40 1 44 0 0 8320 0 47 24 0 0 4
492 350
565 350
565 442
588 442
13 2 45 0 0 4224 0 50 24 0 0 4
895 368
576 368
576 451
588 451
39 3 31 0 0 8320 0 47 24 0 0 4
492 359
554 359
554 460
588 460
44 17 46 0 0 12416 0 47 50 0 0 4
492 314
615 314
615 404
895 404
61 3 47 0 0 8320 0 47 22 0 0 6
336 239
336 234
72 234
72 498
127 498
127 517
1 33 48 0 0 12416 0 58 47 0 0 5
600 614
600 615
523 615
523 413
492 413
1 34 49 0 0 8320 0 57 47 0 0 4
598 586
533 586
533 404
492 404
2 0 5 0 0 0 0 36 0 0 74 2
726 614
735 614
2 1 5 0 0 0 0 38 37 0 0 3
726 586
735 586
735 626
1 0 50 0 0 4096 0 60 0 0 77 2
656 576
656 586
1 0 51 0 0 4096 0 59 0 0 78 2
672 577
672 614
1 2 50 0 0 4224 0 38 57 0 0 2
692 586
634 586
1 2 51 0 0 4224 0 36 58 0 0 2
692 614
636 614
0 2 4 0 0 0 0 0 59 80 0 3
664 532
672 532
672 541
1 2 4 0 0 0 0 8 60 0 0 4
664 525
664 532
656 532
656 540
58 1 52 0 0 4224 0 47 34 0 0 3
363 239
363 205
346 205
57 1 53 0 0 4224 0 47 33 0 0 3
372 239
372 175
345 175
2 2 54 0 0 4224 0 34 56 0 0 4
326 205
331 205
331 205
326 205
2 2 55 0 0 12416 0 55 33 0 0 4
326 175
331 175
331 175
325 175
1 0 5 0 0 0 0 56 0 0 86 2
290 205
281 205
1 1 5 0 0 0 0 55 35 0 0 3
290 175
281 175
281 207
0 2 4 0 0 0 0 0 54 95 0 2
385 527
385 535
0 1 33 0 0 0 0 0 54 40 0 2
385 578
385 571
9 43 56 0 0 4224 0 50 47 0 0 4
895 332
631 332
631 323
492 323
7 42 57 0 0 4224 0 50 47 0 0 4
895 314
622 314
622 332
492 332
3 0 5 0 0 0 0 31 0 0 92 3
336 579
336 501
369 501
5 0 5 0 0 0 0 29 0 0 93 3
417 502
417 501
369 501
0 1 5 0 0 0 0 0 27 94 0 2
369 470
369 507
25 20 5 0 0 0 0 47 47 0 0 4
390 451
390 470
345 470
345 451
0 2 4 0 0 0 0 0 31 109 0 4
385 480
385 527
345 527
345 579
18 4 58 0 0 4224 0 47 31 0 0 2
327 451
327 579
5 17 59 0 0 4224 0 31 47 0 0 2
318 579
318 451
2 0 3 0 0 0 0 30 0 0 99 3
884 240
884 226
838 226
1 11 3 0 0 4224 0 5 50 0 0 3
838 212
838 350
895 350
1 0 5 0 0 0 0 30 0 0 112 2
884 258
884 269
4 0 3 0 0 0 0 50 0 0 99 2
895 287
838 287
7 0 5 0 0 0 0 48 0 0 42 2
184 377
240 377
21 4 60 0 0 8320 0 47 29 0 0 4
354 451
354 463
426 463
426 502
29 3 61 0 0 12416 0 47 29 0 0 4
426 451
426 458
435 458
435 502
31 2 62 0 0 4224 0 47 29 0 0 2
444 451
444 502
32 1 63 0 0 4224 0 47 29 0 0 2
453 451
453 502
2 56 64 0 0 8320 0 15 47 0 0 3
427 143
390 143
390 239
1 41 5 0 0 0 0 28 47 0 0 3
585 343
585 341
492 341
19 0 4 0 0 0 0 47 0 0 110 3
336 451
336 480
404 480
26 1 4 0 0 0 0 47 11 0 0 5
399 451
399 480
404 480
404 481
409 481
5 6 4 0 0 0 0 48 48 0 0 4
184 395
191 395
191 386
184 386
0 2 5 0 0 0 0 0 50 113 0 3
816 386
816 269
895 269
15 1 5 0 0 0 0 50 25 0 0 3
895 386
816 386
816 461
1 10 2 0 0 0 0 3 50 0 0 2
889 341
895 341
5 8 65 0 0 4224 0 47 48 0 0 4
280 314
185 314
185 368
184 368
6 1 66 0 0 4224 0 47 48 0 0 4
280 323
94 323
94 368
100 368
8 4 67 0 0 12416 0 47 48 0 0 6
280 341
198 341
198 430
84 430
84 395
100 395
4 2 68 0 0 4224 0 47 48 0 0 4
280 305
89 305
89 377
100 377
2 2 4 0 0 0 0 53 52 0 0 4
801 225
801 216
764 216
764 226
1 0 37 0 0 0 0 53 0 0 123 2
801 261
801 296
1 0 30 0 0 4096 0 52 0 0 122 2
764 262
764 277
8 3 30 0 0 16512 0 22 50 0 0 11
172 517
172 497
250 497
250 624
505 624
505 386
654 386
654 277
764 277
764 278
895 278
5 37 37 0 0 4224 0 50 47 0 0 4
895 296
604 296
604 377
492 377
12 55 69 0 0 12416 0 50 47 0 0 5
895 359
744 359
744 164
399 164
399 239
14 54 70 0 0 12416 0 50 47 0 0 5
895 377
737 377
737 169
408 169
408 239
16 53 71 0 0 12416 0 50 47 0 0 5
895 395
731 395
731 176
417 176
417 239
18 52 72 0 0 12416 0 50 47 0 0 5
895 413
726 413
726 182
426 182
426 239
20 51 73 0 0 12416 0 50 47 0 0 5
895 431
719 431
719 188
435 188
435 239
22 50 74 0 0 12416 0 50 47 0 0 5
895 449
712 449
712 194
444 194
444 239
21 49 75 0 0 12416 0 50 47 0 0 5
895 440
705 440
705 202
453 202
453 239
19 46 76 0 0 4224 0 50 47 0 0 4
895 422
595 422
595 296
492 296
64 1 4 0 0 0 0 47 13 0 0 2
382 239
382 148
1 1 5 0 0 0 0 41 40 0 0 2
357 88
357 83
2 0 4 0 0 0 0 40 0 0 135 2
357 65
357 51
1 5 4 0 0 0 0 14 45 0 0 2
373 51
338 51
2 0 34 0 0 0 0 44 0 0 138 2
221 59
221 51
3 0 34 0 0 0 0 45 0 0 138 3
277 83
270 83
270 51
1 2 34 0 0 0 0 45 43 0 0 4
277 51
221 51
221 52
41 52
2 0 5 0 0 0 0 45 0 0 140 4
277 67
256 67
256 87
221 87
1 1 5 0 0 0 0 42 44 0 0 2
221 90
221 77
4
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 38
938 331 1019 415
942 335 1014 399
38 Extension
Flat Flex
Cable
.5mm - 24
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
715 30 754 48
718 33 750 45
5 =1.8V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
655 20 694 38
658 23 690 35
5 =2.5V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
392 33 431 51
395 36 427 48
5 =3.3V
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
