CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 230 10
176 83 1438 857
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
21 1Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
77070354 0
0
2 

2 

0
0
0
19
9 Schottky~
219 170 119 0 2 5
0 3 4
0
0 0 576 90
10 PMEG2015EJ
5 -1 75 7
2 D1
13 -7 27 1
0
0
11 %D %1 %2 %M
0
0
12 SM/D/SC90/KA
5

0 -54 -44 -54 -44 0
68 0 0 0 0 1 0 0
1 D
5690 0 0
2
39610.5 0
0
5 SIP2~
219 54 194 0 2 5
0 13 7
0
0 0 352 180
12 Flap Control
-47 -20 37 -12
4 CON1
-20 -30 8 -22
0
0
0
0
0
5 Pad-2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
3 CON
5617 0 0
2
39610 0
0
10 Capacitor~
219 78 268 0 2 5
0 2 7
0
0 0 832 90
4 22nF
10 1 38 9
2 C2
17 -9 31 -1
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3903 0 0
2
39610 1
0
10 N-EMOS 3T~
219 192 230 0 3 7
0 3 12 2
0
0 0 832 0
9 ZXMN2B01F
11 2 74 10
2 Q1
12 -10 26 -2
31 IC-MOSFET N-ch 20V-2.1A-LogicOn
-110 -48 107 -40
0
17 %D %1 %2 %3 %3 %M
0
0
9 SOT23/GSD
7

0 -51 -48 -36 -51 -48 -36 0
77 0 0 0 1 1 0 0
1 Q
4452 0 0
2
39610 2
0
7 Ground~
168 145 307 0 1 3
0 2
0
0 0 53344 512
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6282 0 0
2
39610 3
0
5 SIP2~
219 230 87 0 2 5
0 4 3
0
0 0 352 0
14 Flapping Motor
-49 -22 49 -14
4 CON2
-14 -20 14 -12
0
0
0
0
0
5 Pad-2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
3 CON
7187 0 0
2
39610 4
0
7 Ground~
168 304 59 0 1 3
0 2
0
0 0 53344 512
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6866 0 0
2
39610 5
0
5 SIP2~
219 303 38 0 2 5
0 2 4
0
0 0 864 602
5 <4.2V
-21 -19 14 -11
7 Battery
-28 -29 21 -21
0
0
0
0
0
5 Pad-2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
3 CON
7670 0 0
2
39610 6
0
10 Capacitor~
219 130 118 0 2 5
0 3 4
0
0 0 832 90
3 1nF
11 0 32 8
2 C1
15 -9 29 -1
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
951 0 0
2
39610 7
0
5 SIP2~
219 454 82 0 2 5
0 9 8
0
0 0 352 692
14 Steering Motor
-48 -22 50 -14
4 CON4
-14 -20 14 -12
0
0
0
0
0
5 Pad-2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
3 CON
9536 0 0
2
39610 9
0
5 SIP2~
219 256 197 0 2 5
0 11 10
0
0 0 352 180
13 Steer Control
-46 -20 45 -12
4 CON3
-20 -30 8 -22
0
0
0
0
0
5 Pad-2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
3 CON
5495 0 0
2
39610 10
0
7 Ground~
168 303 304 0 1 3
0 2
0
0 0 53344 512
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8152 0 0
2
39610 11
0
8 H-bridge
94 359 274 0 8 17
0 5 2 6 5 9 4 8 6
8 H-bridge
1 0 4864 0
11 ZXMHC3A01T8
-34 21 43 29
2 H1
-6 -38 8 -30
63 Complementary 30V-2.3A-LogicOn Enhancement Mode MOSFET H-bridge
-220 -57 221 -49
0
0
0
0
4 SM-8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
1 H
6223 0 0
2
39610 12
0
10 Capacitor~
219 427 156 0 2 5
0 9 8
0
0 0 832 180
3 1nF
-11 -18 10 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
9 SM/C/0402
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5441 0 0
2
39610 13
0
9 Resistor~
219 143 191 0 2 5
0 7 3
0
0 0 864 0
3 300
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3189 0 0
2
39610 14
0
9 Resistor~
219 118 239 0 2 5
0 13 12
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8460 0 0
2
39610 15
0
9 Resistor~
219 145 268 0 3 5
0 2 12 -1
0
0 0 864 90
4 100k
4 0 32 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5179 0 0
2
39610 16
0
9 Resistor~
219 289 256 0 2 5
0 11 5
0
0 0 864 0
2 1k
-5 -12 9 -4
2 R4
-5 -23 9 -15
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3593 0 0
2
39610 17
0
9 Resistor~
219 294 226 0 2 5
0 10 6
0
0 0 864 0
2 1k
-8 -12 6 -4
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
9 SM/R/0402
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3928 0 0
2
39610 18
0
28
1 0 3 0 0 4096 0 1 0 0 28 2
171 129
171 153
2 0 4 0 0 4096 0 1 0 0 3 2
171 106
171 83
2 0 4 0 0 8192 0 9 0 0 10 3
130 109
130 83
171 83
1 1 2 0 0 4096 0 8 7 0 0 2
304 47
304 53
2 0 5 0 0 4096 0 18 0 0 18 2
307 256
311 256
2 0 6 0 0 4096 0 19 0 0 17 2
312 226
320 226
0 6 4 0 0 12416 0 0 13 10 0 5
283 49
283 137
403 137
403 274
392 274
2 0 7 0 0 4224 0 3 0 0 23 2
78 259
78 191
0 1 2 0 0 4224 0 0 3 27 0 3
145 293
78 293
78 277
2 1 4 0 0 16 0 8 6 0 0 5
295 47
295 49
171 49
171 83
218 83
2 0 8 0 0 4096 0 14 0 0 13 2
418 156
411 156
0 1 9 0 0 4096 0 0 14 14 0 4
442 156
430 156
430 156
436 156
2 7 8 0 0 8320 0 10 13 0 0 4
442 79
411 79
411 265
392 265
1 5 9 0 0 4224 0 10 13 0 0 3
442 88
442 283
392 283
2 1 10 0 0 8320 0 11 19 0 0 4
260 194
274 194
274 226
276 226
1 1 11 0 0 8320 0 11 18 0 0 4
260 203
266 203
266 256
271 256
3 8 6 0 0 12416 0 13 13 0 0 6
326 274
320 274
320 226
396 226
396 256
392 256
4 1 5 0 0 8320 0 13 13 0 0 4
326 283
311 283
311 256
326 256
2 1 2 0 0 0 0 13 12 0 0 3
326 265
303 265
303 298
2 0 3 0 0 4096 0 15 0 0 25 2
161 191
198 191
0 2 12 0 0 4096 0 0 17 22 0 2
145 239
145 250
2 2 12 0 0 4224 0 4 16 0 0 2
174 239
136 239
2 1 7 0 0 0 0 2 15 0 0 2
58 191
125 191
1 1 13 0 0 8320 0 16 2 0 0 4
100 239
90 239
90 200
58 200
1 2 3 0 0 4224 0 4 6 0 0 3
198 212
198 92
218 92
1 0 2 0 0 0 0 5 0 0 27 2
145 301
145 293
1 3 2 0 0 0 0 17 4 0 0 4
145 286
145 293
198 293
198 248
1 0 3 0 0 0 0 9 0 0 25 3
130 127
130 153
198 153
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
